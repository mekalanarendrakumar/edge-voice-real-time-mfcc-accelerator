// Wake Word RTL placeholder
module wake_word();
// ...implementation...
endmodule
